library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.ReedSolomon.all;

-- Inversion table used by the Chien Search and Forney's algorithm module

-- output = (input)^-1

entity inversion_table is
  port (
    input  : in  field_element;
    output : out field_element);
end inversion_table;

architecture inversion_table of inversion_table is
  type rom_table is array (0 to N_LENGTH) of field_element;
  constant inversion : rom_table := ("00000000",
                                     "00000001",
                                     "10001110",
                                     "11110100",
                                     "01000111",
                                     "10100111",
                                     "01111010",
                                     "10111010",
                                     "10101101",
                                     "10011101",
                                     "11011101",
                                     "10011000",
                                     "00111101",
                                     "10101010",
                                     "01011101",
                                     "10010110",
                                     "11011000",
                                     "01110010",
                                     "11000000",
                                     "01011000",
                                     "11100000",
                                     "00111110",
                                     "01001100",
                                     "01100110",
                                     "10010000",
                                     "11011110",
                                     "01010101",
                                     "10000000",
                                     "10100000",
                                     "10000011",
                                     "01001011",
                                     "00101010",
                                     "01101100",
                                     "11101101",
                                     "00111001",
                                     "01010001",
                                     "01100000",
                                     "01010110",
                                     "00101100",
                                     "10001010",
                                     "01110000",
                                     "11010000",
                                     "00011111",
                                     "01001010",
                                     "00100110",
                                     "10001011",
                                     "00110011",
                                     "01101110",
                                     "01001000",
                                     "10001001",
                                     "01101111",
                                     "00101110",
                                     "10100100",
                                     "11000011",
                                     "01000000",
                                     "01011110",
                                     "01010000",
                                     "00100010",
                                     "11001111",
                                     "10101001",
                                     "10101011",
                                     "00001100",
                                     "00010101",
                                     "11100001",
                                     "00110110",
                                     "01011111",
                                     "11111000",
                                     "11010101",
                                     "10010010",
                                     "01001110",
                                     "10100110",
                                     "00000100",
                                     "00110000",
                                     "10001000",
                                     "00101011",
                                     "00011110",
                                     "00010110",
                                     "01100111",
                                     "01000101",
                                     "10010011",
                                     "00111000",
                                     "00100011",
                                     "01101000",
                                     "10001100",
                                     "10000001",
                                     "00011010",
                                     "00100101",
                                     "01100001",
                                     "00010011",
                                     "11000001",
                                     "11001011",
                                     "01100011",
                                     "10010111",
                                     "00001110",
                                     "00110111",
                                     "01000001",
                                     "00100100",
                                     "01010111",
                                     "11001010",
                                     "01011011",
                                     "10111001",
                                     "11000100",
                                     "00010111",
                                     "01001101",
                                     "01010010",
                                     "10001101",
                                     "11101111",
                                     "10110011",
                                     "00100000",
                                     "11101100",
                                     "00101111",
                                     "00110010",
                                     "00101000",
                                     "11010001",
                                     "00010001",
                                     "11011001",
                                     "11101001",
                                     "11111011",
                                     "11011010",
                                     "01111001",
                                     "11011011",
                                     "01110111",
                                     "00000110",
                                     "10111011",
                                     "10000100",
                                     "11001101",
                                     "11111110",
                                     "11111100",
                                     "00011011",
                                     "01010100",
                                     "10100001",
                                     "00011101",
                                     "01111100",
                                     "11001100",
                                     "11100100",
                                     "10110000",
                                     "01001001",
                                     "00110001",
                                     "00100111",
                                     "00101101",
                                     "01010011",
                                     "01101001",
                                     "00000010",
                                     "11110101",
                                     "00011000",
                                     "11011111",
                                     "01000100",
                                     "01001111",
                                     "10011011",
                                     "10111100",
                                     "00001111",
                                     "01011100",
                                     "00001011",
                                     "11011100",
                                     "10111101",
                                     "10010100",
                                     "10101100",
                                     "00001001",
                                     "11000111",
                                     "10100010",
                                     "00011100",
                                     "10000010",
                                     "10011111",
                                     "11000110",
                                     "00110100",
                                     "11000010",
                                     "01000110",
                                     "00000101",
                                     "11001110",
                                     "00111011",
                                     "00001101",
                                     "00111100",
                                     "10011100",
                                     "00001000",
                                     "10111110",
                                     "10110111",
                                     "10000111",
                                     "11100101",
                                     "11101110",
                                     "01101011",
                                     "11101011",
                                     "11110010",
                                     "10111111",
                                     "10101111",
                                     "11000101",
                                     "01100100",
                                     "00000111",
                                     "01111011",
                                     "10010101",
                                     "10011010",
                                     "10101110",
                                     "10110110",
                                     "00010010",
                                     "01011001",
                                     "10100101",
                                     "00110101",
                                     "01100101",
                                     "10111000",
                                     "10100011",
                                     "10011110",
                                     "11010010",
                                     "11110111",
                                     "01100010",
                                     "01011010",
                                     "10000101",
                                     "01111101",
                                     "10101000",
                                     "00111010",
                                     "00101001",
                                     "01110001",
                                     "11001000",
                                     "11110110",
                                     "11111001",
                                     "01000011",
                                     "11010111",
                                     "11010110",
                                     "00010000",
                                     "01110011",
                                     "01110110",
                                     "01111000",
                                     "10011001",
                                     "00001010",
                                     "00011001",
                                     "10010001",
                                     "00010100",
                                     "00111111",
                                     "11100110",
                                     "11110000",
                                     "10000110",
                                     "10110001",
                                     "11100010",
                                     "11110001",
                                     "11111010",
                                     "01110100",
                                     "11110011",
                                     "10110100",
                                     "01101101",
                                     "00100001",
                                     "10110010",
                                     "01101010",
                                     "11100011",
                                     "11100111",
                                     "10110101",
                                     "11101010",
                                     "00000011",
                                     "10001111",
                                     "11010011",
                                     "11001001",
                                     "01000010",
                                     "11010100",
                                     "11101000",
                                     "01110101",
                                     "01111111",
                                     "11111111",
                                     "01111110",
                                     "11111101");

begin
  output <= inversion(to_integer(unsigned(input)));
end inversion_table;
